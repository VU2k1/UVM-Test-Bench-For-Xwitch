`include "uvm_macros.svh"
import xsw_transaction::*;
import uvm_pkg::*;

typedef uvm_sequencer #(transaction) xsw_sequencer;
